module flipflop ( 
	q,
	clock,
	d
	) ;

inout  q;
input  clock;
input  d;
