module comparador ( 
	x,
	y,
	z,
	display
	) ;

input [3:0] x;
input [3:0] y;
input [3:0] z;
inout [6:0] display;
