module compuertas ( 
	a,
	yand,
	yor,
	ynand,
	ynor,
	yxor,
	yxnor
	) ;

input [3:0] a;
inout  yand;
inout  yor;
inout  ynand;
inout  ynor;
inout  yxor;
inout  yxnor;
