module compuertas ( 
	a,
	b,
	c,
	d,
	andx,
	orx,
	nandx,
	norx,
	xorx,
	xnorx
	) ;

input  a;
input  b;
input  c;
input  d;
inout  andx;
inout  orx;
inout  nandx;
inout  norx;
inout  xorx;
inout  xnorx;
