
--  CYPRESS NOVA XVL Structural Architecture

--  JED2VHD Reverse Assembler - 6.3 IR 35


--    VHDL File: Sumador completo.vhd

--    Date: Wed Nov 10 02:52:01 2021

--  Disassembly from Jedec file for: c22v10

--  Device Ordercode is: PALC22V10D-25PC
library ieee;
use ieee.std_logic_1164.all;

library primitive;
use primitive.primitive.all;


-- Beginning Test Bench Header

ENTITY suma IS
    PORT (
	                  a3 :    in std_logic ;
	                  a2 :    in std_logic ;
	                  a1 :    in std_logic ;
	                  a0 :    in std_logic ;
	                  b3 :    in std_logic ;
	                  b2 :    in std_logic ;
	                  b1 :    in std_logic ;
	                  b0 :    in std_logic ;
	                 cin :    in std_logic ;
	                  s0 : inout std_logic ;
	                  s1 : inout std_logic ;
	                  s2 : inout std_logic ;
	                  s3 : inout std_logic ;
	               cout0 : inout std_logic ;
	               cout2 : inout std_logic ;
	               cout3 : inout std_logic
    );
END suma;

-- End of Test Bench Header

ARCHITECTURE DSMB of suma is

	signal jed_node1	: std_logic:='0' ; -- b3
	signal jed_node2	: std_logic:='0' ; -- b2
	signal jed_node3	: std_logic:='0' ; -- a3
	signal jed_node4	: std_logic:='0' ; -- a2
	signal jed_node5	: std_logic:='0' ; -- b1
	signal jed_node6	: std_logic:='0' ; -- b0
	signal jed_node7	: std_logic:='0' ; -- a1
	signal jed_node8	: std_logic:='0' ; -- a0
	signal jed_node9	: std_logic:='0' ;
	signal jed_node10	: std_logic:='0' ;
	signal jed_node11	: std_logic:='0' ;
	signal jed_node12	: std_logic:='0' ;
	signal jed_node13	: std_logic:='0' ;
	signal jed_node18	: std_logic:='0' ;
	signal jed_node19	: std_logic:='0' ;
	signal jed_node23	: std_logic:='0' ; -- cin
	signal jed_node24	: std_logic:='0' ;

	for all: c22v10m use entity primitive.c22v10m (sim);

SIGNAL  one:std_logic:='1';
SIGNAL  zero:std_logic:='0';
SIGNAL  jed_oept_1:std_logic:='0';
--Attribute PIN_NUMBERS of b3:SIGNAL is "0001";

SIGNAL  jed_oept_2:std_logic:='0';
--Attribute PIN_NUMBERS of b2:SIGNAL is "0002";

SIGNAL  jed_oept_3:std_logic:='0';
--Attribute PIN_NUMBERS of a3:SIGNAL is "0003";

SIGNAL  jed_oept_4:std_logic:='0';
--Attribute PIN_NUMBERS of a2:SIGNAL is "0004";

SIGNAL  jed_oept_5:std_logic:='0';
--Attribute PIN_NUMBERS of b1:SIGNAL is "0005";

SIGNAL  jed_oept_6:std_logic:='0';
--Attribute PIN_NUMBERS of b0:SIGNAL is "0006";

SIGNAL  jed_oept_7:std_logic:='0';
--Attribute PIN_NUMBERS of a1:SIGNAL is "0007";

SIGNAL  jed_oept_8:std_logic:='0';
--Attribute PIN_NUMBERS of a0:SIGNAL is "0008";

SIGNAL  jed_oept_14:std_logic:='0';
SIGNAL  jed_sum_14,jed_fb_14:std_logic:='0';
--Attribute PIN_NUMBERS of cout3:SIGNAL is "0014";

SIGNAL  jed_oept_15:std_logic:='0';
SIGNAL  jed_sum_15,jed_fb_15:std_logic:='0';
--Attribute PIN_NUMBERS of s2:SIGNAL is "0015";

SIGNAL  jed_oept_16:std_logic:='0';
SIGNAL  jed_sum_16,jed_fb_16:std_logic:='0';
--Attribute PIN_NUMBERS of s3:SIGNAL is "0016";

SIGNAL  jed_oept_17:std_logic:='0';
SIGNAL  jed_sum_17,jed_fb_17:std_logic:='0';
--Attribute PIN_NUMBERS of cout2:SIGNAL is "0017";

SIGNAL  jed_oept_20:std_logic:='0';
SIGNAL  jed_sum_20,jed_fb_20:std_logic:='0';
--Attribute PIN_NUMBERS of cout0:SIGNAL is "0020";

SIGNAL  jed_oept_21:std_logic:='0';
SIGNAL  jed_sum_21,jed_fb_21:std_logic:='0';
--Attribute PIN_NUMBERS of s1:SIGNAL is "0021";

SIGNAL  jed_oept_22:std_logic:='0';
SIGNAL  jed_sum_22,jed_fb_22:std_logic:='0';
--Attribute PIN_NUMBERS of s0:SIGNAL is "0022";

SIGNAL  jed_oept_23:std_logic:='0';
SIGNAL  jed_sum_23,jed_fb_23:std_logic:='0';
--Attribute PIN_NUMBERS of cin:SIGNAL is "0023";

SIGNAL  jed_oept_25:std_logic:='0';
SIGNAL  jed_node25,jed_sum_25:std_logic:='0';
SIGNAL  jed_oept_26:std_logic:='0';
SIGNAL  jed_node26,jed_sum_26:std_logic:='0';

BEGIN
jed_node1 <= b3 ;
jed_node2 <= b2 ;
jed_node3 <= a3 ;
jed_node4 <= a2 ;
jed_node5 <= b1 ;
jed_node6 <= b0 ;
jed_node7 <= a1 ;
jed_node8 <= a0 ;
jed_node23 <= cin ;
Mcell_14:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_14,
     clk=>jed_node1,
     oe=>jed_oept_14,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>cout3,
     fb=>jed_fb_14
   );

Mcell_15:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_15,
     clk=>jed_node1,
     oe=>jed_oept_15,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>s2,
     fb=>jed_fb_15
   );

Mcell_16:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_16,
     clk=>jed_node1,
     oe=>jed_oept_16,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>s3,
     fb=>jed_fb_16
   );

Mcell_17:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_17,
     clk=>jed_node1,
     oe=>jed_oept_17,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>cout2,
     fb=>jed_fb_17
   );

Mcell_20:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_20,
     clk=>jed_node1,
     oe=>jed_oept_20,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>cout0,
     fb=>jed_fb_20
   );

Mcell_21:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_21,
     clk=>jed_node1,
     oe=>jed_oept_21,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>s1,
     fb=>jed_fb_21
   );

Mcell_22:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_22,
     clk=>jed_node1,
     oe=>jed_oept_22,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>s0,
     fb=>jed_fb_22
   );

Mcell_23:c22v10m
generic map(comb,
   ninv,
   xpin,
   	25 ns, --tpd
	25 ns, --tea
	25 ns, --ter
	15 ns, --tco
	18 ns, --ts
	0 ns, --th
	14 ns, --twh
	14 ns, --twl
	13 ns, --tcf
	25 ns, --taw
	25 ns, --tar
	25 ns, --tap
	25 ns  --tspr
)
port map(
     d=>jed_sum_23,
     clk=>jed_node1,
     oe=>jed_oept_23,
     ss=>jed_sum_26,
     ar=>jed_sum_25,
     y=>jed_node23,
     fb=>jed_fb_23
   );

jed_node25<=jed_sum_25;
jed_node26<=jed_sum_26;
jed_oept_14<=(one);

jed_sum_14<= (((jed_node1) and (jed_fb_23) and (jed_node2)) or
((jed_fb_23) and (jed_node2) and (jed_node3)) or
((jed_node1) and (jed_fb_23) and (jed_node4)) or
((jed_node1) and (jed_node2) and (jed_node4)) or
((jed_fb_23) and (jed_node3) and (jed_node4)) or
((jed_node2) and (jed_node3) and (jed_node4)) or
((jed_node1) and (jed_node3)));

jed_oept_15<=(one);

jed_sum_15<= (((jed_fb_23) and (jed_node2) and (jed_node4)) or
((jed_fb_23) and not(jed_node2) and not(jed_node4)) or
(not(jed_fb_23) and (jed_node2) and not(jed_node4)) or
(not(jed_fb_23) and not(jed_node2) and (jed_node4)));

jed_oept_16<=(one);

jed_sum_16<= (((jed_node1) and (jed_fb_23) and (jed_node2) and (jed_node3)
) or
((jed_node1) and (jed_fb_23) and (jed_node3) and (jed_node4)
) or
((jed_node1) and (jed_node2) and (jed_node3) and (jed_node4)
) or
((jed_node1) and not(jed_node2) and not(jed_node3) and not(jed_node4)
) or
(not(jed_node1) and (jed_fb_23) and (jed_node2) and not(jed_node3)
) or
(not(jed_node1) and (jed_fb_23) and not(jed_node3) and (jed_node4)
) or
(not(jed_node1) and (jed_node2) and not(jed_node3) and (jed_node4)
) or
(not(jed_node1) and not(jed_node2) and (jed_node3) and not(jed_node4)
) or
((jed_node1) and not(jed_fb_23) and not(jed_node3) and not(jed_node4)
) or
((jed_node1) and not(jed_fb_23) and not(jed_node2) and not(jed_node3)
) or
(not(jed_node1) and not(jed_fb_23) and (jed_node3) and not(jed_node4)
) or
(not(jed_node1) and not(jed_fb_23) and not(jed_node2)
 and (jed_node3)));

jed_oept_17<=(one);

jed_sum_17<= (((jed_fb_23) and (jed_node2)) or
((jed_fb_23) and (jed_node4)) or
((jed_node2) and (jed_node4)));

jed_oept_20<=(one);

jed_sum_20<= (((jed_fb_23) and (jed_node6)) or
((jed_fb_23) and (jed_node8)) or
((jed_node6) and (jed_node8)));

jed_oept_21<=(one);

jed_sum_21<= (((jed_fb_23) and (jed_node5) and (jed_node6) and (jed_node7)
) or
((jed_fb_23) and (jed_node5) and (jed_node7) and (jed_node8)
) or
((jed_node5) and (jed_node6) and (jed_node7) and (jed_node8)
) or
((jed_node5) and not(jed_node6) and not(jed_node7) and not(jed_node8)
) or
((jed_fb_23) and not(jed_node5) and (jed_node6) and not(jed_node7)
) or
((jed_fb_23) and not(jed_node5) and not(jed_node7) and (jed_node8)
) or
(not(jed_node5) and (jed_node6) and not(jed_node7) and (jed_node8)
) or
(not(jed_node5) and not(jed_node6) and (jed_node7) and not(jed_node8)
) or
(not(jed_fb_23) and (jed_node5) and not(jed_node7) and not(jed_node8)
) or
(not(jed_fb_23) and (jed_node5) and not(jed_node6) and not(jed_node7)
) or
(not(jed_fb_23) and not(jed_node5) and (jed_node7) and not(jed_node8)
) or
(not(jed_fb_23) and not(jed_node5) and not(jed_node6)
 and (jed_node7)));

jed_oept_22<=(one);

jed_sum_22<= (((jed_fb_23) and (jed_node6) and (jed_node8)) or
((jed_fb_23) and not(jed_node6) and not(jed_node8)) or
(not(jed_fb_23) and (jed_node6) and not(jed_node8)) or
(not(jed_fb_23) and not(jed_node6) and (jed_node8)));

jed_oept_23<=(one);

jed_sum_23<= (((jed_fb_23) and (jed_node5) and (jed_node6)) or
((jed_fb_23) and (jed_node6) and (jed_node7)) or
((jed_fb_23) and (jed_node5) and (jed_node8)) or
((jed_node5) and (jed_node6) and (jed_node8)) or
((jed_fb_23) and (jed_node7) and (jed_node8)) or
((jed_node6) and (jed_node7) and (jed_node8)) or
((jed_node5) and (jed_node7)));

end DSMB;
