module rs_ff ( 
	clk,
	r,
	s,
	q,
	qnot
	) ;

input  clk;
input  r;
input  s;
inout  q;
inout  qnot;
