module comparador ( 
	x,
	y,
	mayor,
	menor,
	igual,
	display
	) ;

input [3:0] x;
input [3:0] y;
inout  mayor;
inout  menor;
inout  igual;
inout [6:0] display;
