module resta ( 
	a,
	b,
	resta,
	carry
	) ;

input  a;
input  b;
inout  resta;
inout  carry;
