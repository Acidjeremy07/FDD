module suma ( 
	a0,
	a1,
	a2,
	a3,
	b0,
	b1,
	b2,
	b3,
	cin0,
	cin1,
	cin2,
	cout0,
	cout1,
	cout2,
	cout3,
	s0,
	s1,
	s2,
	s3
	) ;

input  a0;
input  a1;
input  a2;
input  a3;
input  b0;
input  b1;
input  b2;
input  b3;
input  cin0;
input  cin1;
input  cin2;
inout  cout0;
inout  cout1;
inout  cout2;
inout  cout3;
inout  s0;
inout  s1;
inout  s2;
inout  s3;
