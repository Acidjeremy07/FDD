module multiplexor ( 
	w0,
	w1,
	w2,
	w3,
	selec,
	f
	) ;

input  w0;
input  w1;
input  w2;
input  w3;
input [1:0] selec;
inout  f;
