module compuerta_or ( 
	a,
	b,
	c,
	d,
	salida
	) ;

input  a;
input  b;
input  c;
input  d;
inout  salida;
