module flipflopsrs ( 
	clk,
	rst,
	s,
	r,
	q
	) ;

input  clk;
input  rst;
input  s;
input  r;
inout  q;
