module suma ( 
	a,
	b,
	cin,
	suma,
	carry
	) ;

input  a;
input  b;
input  cin;
inout  suma;
inout  carry;
