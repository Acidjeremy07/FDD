module ffjk ( 
	clk,
	rst,
	j,
	k,
	q
	) ;

input  clk;
input  rst;
input  j;
input  k;
inout  q;
