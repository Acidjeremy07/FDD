module deco ( 
	a,
	b,
	c,
	d,
	e,
	f,
	g,
	x3,
	x2,
	x1,
	x0
	) ;

inout  a;
inout  b;
inout  c;
inout  d;
inout  e;
inout  f;
inout  g;
input  x3;
input  x2;
input  x1;
input  x0;
