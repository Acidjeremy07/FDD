module sr_ff ( 
	s,
	r,
	clock,
	q,
	qbar
	) ;

input  s;
input  r;
input  clock;
inout  q;
inout  qbar;
