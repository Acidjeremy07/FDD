module fft ( 
	t,
	clock,
	q
	) ;

input  t;
input  clock;
inout  q;
