module suma ( 
	a3,
	a2,
	a1,
	a0,
	b3,
	b2,
	b1,
	b0,
	cin,
	s0,
	s1,
	s2,
	s3,
	cout0,
	cout2,
	cout3
	) ;

input  a3;
input  a2;
input  a1;
input  a0;
input  b3;
input  b2;
input  b1;
input  b0;
input  cin;
inout  s0;
inout  s1;
inout  s2;
inout  s3;
inout  cout0;
inout  cout2;
inout  cout3;
