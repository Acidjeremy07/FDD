module mult ( 
	a0,
	a1,
	b0,
	b1,
	p0,
	p1,
	p2,
	p3
	) ;

input  a0;
input  a1;
input  b0;
input  b1;
inout  p0;
inout  p1;
inout  p2;
inout  p3;
