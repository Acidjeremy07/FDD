module flipflop ( 
	q,
	clk,
	rst,
	d
	) ;

inout  q;
input  clk;
input  rst;
input  d;
