module compuerta_xor ( 
	a,
	b,
	c,
	d,
	salida
	) ;

input  a;
input  b;
input  c;
input  d;
inout  salida;
