module suma ( 
	x,
	y,
	s,
	a
	) ;

input  x;
input  y;
inout  s;
inout  a;
