module resta ( 
	resta,
	cout,
	a,
	b,
	cin
	) ;

inout  resta;
inout  cout;
input  a;
input  b;
input  cin;
